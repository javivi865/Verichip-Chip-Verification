module verichip4_binds;

bind verichip4 verichip4_cov verichip4_cov (.*);

endmodule
